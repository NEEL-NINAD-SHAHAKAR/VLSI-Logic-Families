magic
tech scmos
timestamp 1663573099
<< error_s >>
rect 6 20 13 21
rect 18 20 22 21
rect 23 18 24 31
rect 43 20 50 21
rect 51 18 52 31
rect 60 18 61 31
rect 62 20 69 21
rect 71 20 78 21
rect 79 18 80 31
rect 88 18 89 31
rect 90 20 97 21
rect 99 20 106 21
rect 107 18 108 31
rect 116 18 117 31
rect 118 20 125 21
rect 127 20 134 21
<< error_ps >>
rect 15 20 18 21
rect 32 18 33 31
rect 34 20 41 21
<< metal1 >>
rect -4 14 4 18
rect 136 14 144 18
use CMOS_INV  CMOS_INV_0
array 0 4 28 0 0 37
timestamp 1663501662
transform 1 0 4 0 1 18
box -4 -18 24 19
<< labels >>
rlabel space 70 35 70 35 5 SRC
rlabel space 70 2 70 2 1 GND
rlabel metal1 -2 16 -2 16 3 X
rlabel metal1 142 16 142 16 7 Y
<< end >>
