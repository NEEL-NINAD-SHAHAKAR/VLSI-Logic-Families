magic
tech scmos
timestamp 1664280382
<< nwell >>
rect -22 3 30 34
<< polysilicon >>
rect -5 25 -3 27
rect 9 25 11 27
rect -5 -9 -3 9
rect 9 -9 11 9
rect -5 -28 -3 -25
rect 9 -28 11 -25
<< ndiffusion >>
rect -22 -15 -5 -9
rect -22 -19 -12 -15
rect -8 -19 -5 -15
rect -22 -25 -5 -19
rect -3 -20 9 -9
rect -3 -24 1 -20
rect 5 -24 9 -20
rect -3 -25 9 -24
rect 11 -15 30 -9
rect 11 -19 14 -15
rect 18 -19 30 -15
rect 11 -25 30 -19
<< pdiffusion >>
rect -22 18 -5 25
rect -22 14 -12 18
rect -8 14 -5 18
rect -22 9 -5 14
rect -3 9 9 25
rect 11 18 30 25
rect 11 14 14 18
rect 18 14 30 18
rect 11 9 30 14
<< metal1 >>
rect -22 35 30 40
rect -12 33 -8 35
rect -12 18 -8 29
rect 14 3 18 14
rect -22 -1 -9 3
rect 1 -1 30 3
rect 1 -4 5 -1
rect -12 -8 5 -4
rect 15 -8 30 -4
rect -12 -15 -8 -8
rect 1 -11 5 -8
rect 1 -15 18 -11
rect 1 -30 5 -24
rect -22 -34 1 -30
rect 5 -34 30 -30
rect -22 -35 30 -34
<< ntransistor >>
rect -5 -25 -3 -9
rect 9 -25 11 -9
<< ptransistor >>
rect -5 9 -3 25
rect 9 9 11 25
<< polycontact >>
rect -9 -1 -5 3
rect 11 -8 15 -4
<< ndcontact >>
rect -12 -19 -8 -15
rect 1 -24 5 -20
rect 14 -19 18 -15
<< pdcontact >>
rect -12 14 -8 18
rect 14 14 18 18
<< psubstratepcontact >>
rect 1 -34 5 -30
<< nsubstratencontact >>
rect -12 29 -8 33
<< labels >>
rlabel metal1 3 37 3 37 5 Vdd
rlabel metal1 -20 1 -20 1 3 A
rlabel metal1 28 -6 28 -6 7 B
rlabel metal1 28 1 28 1 7 Out
rlabel psubstratepcontact 3 -32 3 -32 1 Gnd
<< end >>
