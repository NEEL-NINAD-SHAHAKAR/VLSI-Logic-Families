magic
tech scmos
timestamp 1664793188
<< nwell >>
rect -9 2 28 24
<< polysilicon >>
rect -1 15 1 17
rect 9 15 11 17
rect 19 15 21 17
rect -1 -27 1 4
rect 9 -27 11 4
rect 19 -27 21 4
rect -1 -44 1 -42
rect 9 -44 11 -42
rect 19 -44 21 -42
<< ndiffusion >>
rect -9 -35 -1 -27
rect -9 -39 -7 -35
rect -3 -39 -1 -35
rect -9 -42 -1 -39
rect 1 -42 9 -27
rect 11 -42 19 -27
rect 21 -35 28 -27
rect 21 -39 23 -35
rect 27 -39 28 -35
rect 21 -42 28 -39
<< pdiffusion >>
rect -9 10 -1 15
rect -9 6 -7 10
rect -3 6 -1 10
rect -9 4 -1 6
rect 1 10 9 15
rect 1 6 3 10
rect 7 6 9 10
rect 1 4 9 6
rect 11 10 19 15
rect 11 6 13 10
rect 17 6 19 10
rect 11 4 19 6
rect 21 10 28 15
rect 21 6 23 10
rect 27 6 28 10
rect 21 4 28 6
<< metal1 >>
rect -9 19 3 23
rect 7 19 28 23
rect 3 10 7 19
rect 23 10 27 19
rect -7 1 -3 6
rect 13 1 17 6
rect -7 -3 28 1
rect -9 -10 -5 -6
rect -9 -17 5 -13
rect 13 -35 17 -3
rect -3 -39 17 -35
rect 23 -46 27 -39
rect -9 -50 23 -46
rect 27 -50 28 -46
<< metal2 >>
rect -9 -25 21 -21
<< ntransistor >>
rect -1 -42 1 -27
rect 9 -42 11 -27
rect 19 -42 21 -27
<< ptransistor >>
rect -1 4 1 15
rect 9 4 11 15
rect 19 4 21 15
<< polycontact >>
rect -5 -10 -1 -6
rect 5 -17 9 -13
rect 21 -25 25 -21
<< ndcontact >>
rect -7 -39 -3 -35
rect 23 -39 27 -35
<< pdcontact >>
rect -7 6 -3 10
rect 3 6 7 10
rect 13 6 17 10
rect 23 6 27 10
<< psubstratepcontact >>
rect 23 -50 27 -46
<< nsubstratencontact >>
rect 3 19 7 23
<< labels >>
rlabel metal1 10 21 10 21 5 Vdd
rlabel metal1 10 -48 10 -48 1 Gnd
rlabel metal1 26 -1 26 -1 7 Out
rlabel metal1 -6 -8 -6 -8 3 A
rlabel metal1 -6 -15 -6 -15 3 B
rlabel metal2 -6 -23 -6 -23 3 C
<< end >>
